module sink_32 (
    input logic[31:0] sink_in
); 
endmodule
