module sink_1 (
    input logic [0:0] sink_in
); 
endmodule
