`define GLC_TEST_R 'h0
`define GLC_TEST_R_LSB 0
`define GLC_TEST_R_MSB 31
`define GLC_TEST_VALUE_F_LSB 0
`define GLC_TEST_VALUE_F_MSB 31
`define GLC_GLOBAL_RESET_R 'h4
`define GLC_GLOBAL_RESET_R_LSB 0
`define GLC_GLOBAL_RESET_R_MSB 31
`define GLC_GLOBAL_RESET_CNT_F_LSB 0
`define GLC_GLOBAL_RESET_CNT_F_MSB 31
`define GLC_CGRA_STALL_R 'h8
`define GLC_CGRA_STALL_R_LSB 0
`define GLC_CGRA_STALL_R_MSB 31
`define GLC_CGRA_STALL_STALL_F_LSB 0
`define GLC_CGRA_STALL_STALL_F_MSB 31
`define GLC_GLB_CLK_EN_MASTER_R 'hc
`define GLC_GLB_CLK_EN_MASTER_R_LSB 0
`define GLC_GLB_CLK_EN_MASTER_R_MSB 15
`define GLC_GLB_CLK_EN_MASTER_CLK_EN_F_LSB 0
`define GLC_GLB_CLK_EN_MASTER_CLK_EN_F_MSB 15
`define GLC_GLB_CLK_EN_BANK_MASTER_R 'h10
`define GLC_GLB_CLK_EN_BANK_MASTER_R_LSB 0
`define GLC_GLB_CLK_EN_BANK_MASTER_R_MSB 15
`define GLC_GLB_CLK_EN_BANK_MASTER_CLK_EN_F_LSB 0
`define GLC_GLB_CLK_EN_BANK_MASTER_CLK_EN_F_MSB 15
`define GLC_GLB_PCFG_BROADCAST_STALL_R 'h14
`define GLC_GLB_PCFG_BROADCAST_STALL_R_LSB 0
`define GLC_GLB_PCFG_BROADCAST_STALL_R_MSB 15
`define GLC_GLB_PCFG_BROADCAST_STALL_STALL_F_LSB 0
`define GLC_GLB_PCFG_BROADCAST_STALL_STALL_F_MSB 15
`define GLC_STREAM_START_PULSE_R 'h18
`define GLC_STREAM_START_PULSE_R_LSB 0
`define GLC_STREAM_START_PULSE_R_MSB 31
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_0_F_LSB 0
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_0_F_MSB 0
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_1_F_LSB 1
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_1_F_MSB 1
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_2_F_LSB 2
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_2_F_MSB 2
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_3_F_LSB 3
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_3_F_MSB 3
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_4_F_LSB 4
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_4_F_MSB 4
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_5_F_LSB 5
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_5_F_MSB 5
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_6_F_LSB 6
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_6_F_MSB 6
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_7_F_LSB 7
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_7_F_MSB 7
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_8_F_LSB 8
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_8_F_MSB 8
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_9_F_LSB 9
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_9_F_MSB 9
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_10_F_LSB 10
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_10_F_MSB 10
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_11_F_LSB 11
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_11_F_MSB 11
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_12_F_LSB 12
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_12_F_MSB 12
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_13_F_LSB 13
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_13_F_MSB 13
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_14_F_LSB 14
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_14_F_MSB 14
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_15_F_LSB 15
`define GLC_STREAM_START_PULSE_G2F_GLB_TILE_15_F_MSB 15
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_0_F_LSB 16
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_0_F_MSB 16
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_1_F_LSB 17
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_1_F_MSB 17
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_2_F_LSB 18
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_2_F_MSB 18
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_3_F_LSB 19
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_3_F_MSB 19
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_4_F_LSB 20
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_4_F_MSB 20
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_5_F_LSB 21
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_5_F_MSB 21
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_6_F_LSB 22
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_6_F_MSB 22
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_7_F_LSB 23
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_7_F_MSB 23
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_8_F_LSB 24
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_8_F_MSB 24
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_9_F_LSB 25
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_9_F_MSB 25
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_10_F_LSB 26
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_10_F_MSB 26
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_11_F_LSB 27
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_11_F_MSB 27
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_12_F_LSB 28
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_12_F_MSB 28
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_13_F_LSB 29
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_13_F_MSB 29
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_14_F_LSB 30
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_14_F_MSB 30
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_15_F_LSB 31
`define GLC_STREAM_START_PULSE_F2G_GLB_TILE_15_F_MSB 31
`define GLC_PC_START_PULSE_R 'h1c
`define GLC_PC_START_PULSE_R_LSB 0
`define GLC_PC_START_PULSE_R_MSB 15
`define GLC_PC_START_PULSE_GLB_TILE_0_F_LSB 0
`define GLC_PC_START_PULSE_GLB_TILE_0_F_MSB 0
`define GLC_PC_START_PULSE_GLB_TILE_1_F_LSB 1
`define GLC_PC_START_PULSE_GLB_TILE_1_F_MSB 1
`define GLC_PC_START_PULSE_GLB_TILE_2_F_LSB 2
`define GLC_PC_START_PULSE_GLB_TILE_2_F_MSB 2
`define GLC_PC_START_PULSE_GLB_TILE_3_F_LSB 3
`define GLC_PC_START_PULSE_GLB_TILE_3_F_MSB 3
`define GLC_PC_START_PULSE_GLB_TILE_4_F_LSB 4
`define GLC_PC_START_PULSE_GLB_TILE_4_F_MSB 4
`define GLC_PC_START_PULSE_GLB_TILE_5_F_LSB 5
`define GLC_PC_START_PULSE_GLB_TILE_5_F_MSB 5
`define GLC_PC_START_PULSE_GLB_TILE_6_F_LSB 6
`define GLC_PC_START_PULSE_GLB_TILE_6_F_MSB 6
`define GLC_PC_START_PULSE_GLB_TILE_7_F_LSB 7
`define GLC_PC_START_PULSE_GLB_TILE_7_F_MSB 7
`define GLC_PC_START_PULSE_GLB_TILE_8_F_LSB 8
`define GLC_PC_START_PULSE_GLB_TILE_8_F_MSB 8
`define GLC_PC_START_PULSE_GLB_TILE_9_F_LSB 9
`define GLC_PC_START_PULSE_GLB_TILE_9_F_MSB 9
`define GLC_PC_START_PULSE_GLB_TILE_10_F_LSB 10
`define GLC_PC_START_PULSE_GLB_TILE_10_F_MSB 10
`define GLC_PC_START_PULSE_GLB_TILE_11_F_LSB 11
`define GLC_PC_START_PULSE_GLB_TILE_11_F_MSB 11
`define GLC_PC_START_PULSE_GLB_TILE_12_F_LSB 12
`define GLC_PC_START_PULSE_GLB_TILE_12_F_MSB 12
`define GLC_PC_START_PULSE_GLB_TILE_13_F_LSB 13
`define GLC_PC_START_PULSE_GLB_TILE_13_F_MSB 13
`define GLC_PC_START_PULSE_GLB_TILE_14_F_LSB 14
`define GLC_PC_START_PULSE_GLB_TILE_14_F_MSB 14
`define GLC_PC_START_PULSE_GLB_TILE_15_F_LSB 15
`define GLC_PC_START_PULSE_GLB_TILE_15_F_MSB 15
`define GLC_STRM_F2G_IER_R 'h20
`define GLC_STRM_F2G_IER_R_LSB 0
`define GLC_STRM_F2G_IER_R_MSB 15
`define GLC_STRM_F2G_IER_TILE_0_F_LSB 0
`define GLC_STRM_F2G_IER_TILE_0_F_MSB 0
`define GLC_STRM_F2G_IER_TILE_1_F_LSB 1
`define GLC_STRM_F2G_IER_TILE_1_F_MSB 1
`define GLC_STRM_F2G_IER_TILE_2_F_LSB 2
`define GLC_STRM_F2G_IER_TILE_2_F_MSB 2
`define GLC_STRM_F2G_IER_TILE_3_F_LSB 3
`define GLC_STRM_F2G_IER_TILE_3_F_MSB 3
`define GLC_STRM_F2G_IER_TILE_4_F_LSB 4
`define GLC_STRM_F2G_IER_TILE_4_F_MSB 4
`define GLC_STRM_F2G_IER_TILE_5_F_LSB 5
`define GLC_STRM_F2G_IER_TILE_5_F_MSB 5
`define GLC_STRM_F2G_IER_TILE_6_F_LSB 6
`define GLC_STRM_F2G_IER_TILE_6_F_MSB 6
`define GLC_STRM_F2G_IER_TILE_7_F_LSB 7
`define GLC_STRM_F2G_IER_TILE_7_F_MSB 7
`define GLC_STRM_F2G_IER_TILE_8_F_LSB 8
`define GLC_STRM_F2G_IER_TILE_8_F_MSB 8
`define GLC_STRM_F2G_IER_TILE_9_F_LSB 9
`define GLC_STRM_F2G_IER_TILE_9_F_MSB 9
`define GLC_STRM_F2G_IER_TILE_10_F_LSB 10
`define GLC_STRM_F2G_IER_TILE_10_F_MSB 10
`define GLC_STRM_F2G_IER_TILE_11_F_LSB 11
`define GLC_STRM_F2G_IER_TILE_11_F_MSB 11
`define GLC_STRM_F2G_IER_TILE_12_F_LSB 12
`define GLC_STRM_F2G_IER_TILE_12_F_MSB 12
`define GLC_STRM_F2G_IER_TILE_13_F_LSB 13
`define GLC_STRM_F2G_IER_TILE_13_F_MSB 13
`define GLC_STRM_F2G_IER_TILE_14_F_LSB 14
`define GLC_STRM_F2G_IER_TILE_14_F_MSB 14
`define GLC_STRM_F2G_IER_TILE_15_F_LSB 15
`define GLC_STRM_F2G_IER_TILE_15_F_MSB 15
`define GLC_STRM_G2F_IER_R 'h24
`define GLC_STRM_G2F_IER_R_LSB 0
`define GLC_STRM_G2F_IER_R_MSB 15
`define GLC_STRM_G2F_IER_TILE_0_F_LSB 0
`define GLC_STRM_G2F_IER_TILE_0_F_MSB 0
`define GLC_STRM_G2F_IER_TILE_1_F_LSB 1
`define GLC_STRM_G2F_IER_TILE_1_F_MSB 1
`define GLC_STRM_G2F_IER_TILE_2_F_LSB 2
`define GLC_STRM_G2F_IER_TILE_2_F_MSB 2
`define GLC_STRM_G2F_IER_TILE_3_F_LSB 3
`define GLC_STRM_G2F_IER_TILE_3_F_MSB 3
`define GLC_STRM_G2F_IER_TILE_4_F_LSB 4
`define GLC_STRM_G2F_IER_TILE_4_F_MSB 4
`define GLC_STRM_G2F_IER_TILE_5_F_LSB 5
`define GLC_STRM_G2F_IER_TILE_5_F_MSB 5
`define GLC_STRM_G2F_IER_TILE_6_F_LSB 6
`define GLC_STRM_G2F_IER_TILE_6_F_MSB 6
`define GLC_STRM_G2F_IER_TILE_7_F_LSB 7
`define GLC_STRM_G2F_IER_TILE_7_F_MSB 7
`define GLC_STRM_G2F_IER_TILE_8_F_LSB 8
`define GLC_STRM_G2F_IER_TILE_8_F_MSB 8
`define GLC_STRM_G2F_IER_TILE_9_F_LSB 9
`define GLC_STRM_G2F_IER_TILE_9_F_MSB 9
`define GLC_STRM_G2F_IER_TILE_10_F_LSB 10
`define GLC_STRM_G2F_IER_TILE_10_F_MSB 10
`define GLC_STRM_G2F_IER_TILE_11_F_LSB 11
`define GLC_STRM_G2F_IER_TILE_11_F_MSB 11
`define GLC_STRM_G2F_IER_TILE_12_F_LSB 12
`define GLC_STRM_G2F_IER_TILE_12_F_MSB 12
`define GLC_STRM_G2F_IER_TILE_13_F_LSB 13
`define GLC_STRM_G2F_IER_TILE_13_F_MSB 13
`define GLC_STRM_G2F_IER_TILE_14_F_LSB 14
`define GLC_STRM_G2F_IER_TILE_14_F_MSB 14
`define GLC_STRM_G2F_IER_TILE_15_F_LSB 15
`define GLC_STRM_G2F_IER_TILE_15_F_MSB 15
`define GLC_PAR_CFG_G2F_IER_R 'h28
`define GLC_PAR_CFG_G2F_IER_R_LSB 0
`define GLC_PAR_CFG_G2F_IER_R_MSB 15
`define GLC_PAR_CFG_G2F_IER_TILE_0_F_LSB 0
`define GLC_PAR_CFG_G2F_IER_TILE_0_F_MSB 0
`define GLC_PAR_CFG_G2F_IER_TILE_1_F_LSB 1
`define GLC_PAR_CFG_G2F_IER_TILE_1_F_MSB 1
`define GLC_PAR_CFG_G2F_IER_TILE_2_F_LSB 2
`define GLC_PAR_CFG_G2F_IER_TILE_2_F_MSB 2
`define GLC_PAR_CFG_G2F_IER_TILE_3_F_LSB 3
`define GLC_PAR_CFG_G2F_IER_TILE_3_F_MSB 3
`define GLC_PAR_CFG_G2F_IER_TILE_4_F_LSB 4
`define GLC_PAR_CFG_G2F_IER_TILE_4_F_MSB 4
`define GLC_PAR_CFG_G2F_IER_TILE_5_F_LSB 5
`define GLC_PAR_CFG_G2F_IER_TILE_5_F_MSB 5
`define GLC_PAR_CFG_G2F_IER_TILE_6_F_LSB 6
`define GLC_PAR_CFG_G2F_IER_TILE_6_F_MSB 6
`define GLC_PAR_CFG_G2F_IER_TILE_7_F_LSB 7
`define GLC_PAR_CFG_G2F_IER_TILE_7_F_MSB 7
`define GLC_PAR_CFG_G2F_IER_TILE_8_F_LSB 8
`define GLC_PAR_CFG_G2F_IER_TILE_8_F_MSB 8
`define GLC_PAR_CFG_G2F_IER_TILE_9_F_LSB 9
`define GLC_PAR_CFG_G2F_IER_TILE_9_F_MSB 9
`define GLC_PAR_CFG_G2F_IER_TILE_10_F_LSB 10
`define GLC_PAR_CFG_G2F_IER_TILE_10_F_MSB 10
`define GLC_PAR_CFG_G2F_IER_TILE_11_F_LSB 11
`define GLC_PAR_CFG_G2F_IER_TILE_11_F_MSB 11
`define GLC_PAR_CFG_G2F_IER_TILE_12_F_LSB 12
`define GLC_PAR_CFG_G2F_IER_TILE_12_F_MSB 12
`define GLC_PAR_CFG_G2F_IER_TILE_13_F_LSB 13
`define GLC_PAR_CFG_G2F_IER_TILE_13_F_MSB 13
`define GLC_PAR_CFG_G2F_IER_TILE_14_F_LSB 14
`define GLC_PAR_CFG_G2F_IER_TILE_14_F_MSB 14
`define GLC_PAR_CFG_G2F_IER_TILE_15_F_LSB 15
`define GLC_PAR_CFG_G2F_IER_TILE_15_F_MSB 15
`define GLC_GLOBAL_IER_R 'h2c
`define GLC_GLOBAL_IER_R_LSB 0
`define GLC_GLOBAL_IER_R_MSB 2
`define GLC_GLOBAL_IER_STRM_F2G_F_LSB 0
`define GLC_GLOBAL_IER_STRM_F2G_F_MSB 0
`define GLC_GLOBAL_IER_STRM_G2F_F_LSB 1
`define GLC_GLOBAL_IER_STRM_G2F_F_MSB 1
`define GLC_GLOBAL_IER_PAR_CFG_G2F_F_LSB 2
`define GLC_GLOBAL_IER_PAR_CFG_G2F_F_MSB 2
`define GLC_STRM_F2G_ISR_R 'h30
`define GLC_STRM_F2G_ISR_R_LSB 0
`define GLC_STRM_F2G_ISR_R_MSB 15
`define GLC_STRM_F2G_ISR_TILE_0_F_LSB 0
`define GLC_STRM_F2G_ISR_TILE_0_F_MSB 0
`define GLC_STRM_F2G_ISR_TILE_1_F_LSB 1
`define GLC_STRM_F2G_ISR_TILE_1_F_MSB 1
`define GLC_STRM_F2G_ISR_TILE_2_F_LSB 2
`define GLC_STRM_F2G_ISR_TILE_2_F_MSB 2
`define GLC_STRM_F2G_ISR_TILE_3_F_LSB 3
`define GLC_STRM_F2G_ISR_TILE_3_F_MSB 3
`define GLC_STRM_F2G_ISR_TILE_4_F_LSB 4
`define GLC_STRM_F2G_ISR_TILE_4_F_MSB 4
`define GLC_STRM_F2G_ISR_TILE_5_F_LSB 5
`define GLC_STRM_F2G_ISR_TILE_5_F_MSB 5
`define GLC_STRM_F2G_ISR_TILE_6_F_LSB 6
`define GLC_STRM_F2G_ISR_TILE_6_F_MSB 6
`define GLC_STRM_F2G_ISR_TILE_7_F_LSB 7
`define GLC_STRM_F2G_ISR_TILE_7_F_MSB 7
`define GLC_STRM_F2G_ISR_TILE_8_F_LSB 8
`define GLC_STRM_F2G_ISR_TILE_8_F_MSB 8
`define GLC_STRM_F2G_ISR_TILE_9_F_LSB 9
`define GLC_STRM_F2G_ISR_TILE_9_F_MSB 9
`define GLC_STRM_F2G_ISR_TILE_10_F_LSB 10
`define GLC_STRM_F2G_ISR_TILE_10_F_MSB 10
`define GLC_STRM_F2G_ISR_TILE_11_F_LSB 11
`define GLC_STRM_F2G_ISR_TILE_11_F_MSB 11
`define GLC_STRM_F2G_ISR_TILE_12_F_LSB 12
`define GLC_STRM_F2G_ISR_TILE_12_F_MSB 12
`define GLC_STRM_F2G_ISR_TILE_13_F_LSB 13
`define GLC_STRM_F2G_ISR_TILE_13_F_MSB 13
`define GLC_STRM_F2G_ISR_TILE_14_F_LSB 14
`define GLC_STRM_F2G_ISR_TILE_14_F_MSB 14
`define GLC_STRM_F2G_ISR_TILE_15_F_LSB 15
`define GLC_STRM_F2G_ISR_TILE_15_F_MSB 15
`define GLC_STRM_G2F_ISR_R 'h34
`define GLC_STRM_G2F_ISR_R_LSB 0
`define GLC_STRM_G2F_ISR_R_MSB 15
`define GLC_STRM_G2F_ISR_TILE_0_F_LSB 0
`define GLC_STRM_G2F_ISR_TILE_0_F_MSB 0
`define GLC_STRM_G2F_ISR_TILE_1_F_LSB 1
`define GLC_STRM_G2F_ISR_TILE_1_F_MSB 1
`define GLC_STRM_G2F_ISR_TILE_2_F_LSB 2
`define GLC_STRM_G2F_ISR_TILE_2_F_MSB 2
`define GLC_STRM_G2F_ISR_TILE_3_F_LSB 3
`define GLC_STRM_G2F_ISR_TILE_3_F_MSB 3
`define GLC_STRM_G2F_ISR_TILE_4_F_LSB 4
`define GLC_STRM_G2F_ISR_TILE_4_F_MSB 4
`define GLC_STRM_G2F_ISR_TILE_5_F_LSB 5
`define GLC_STRM_G2F_ISR_TILE_5_F_MSB 5
`define GLC_STRM_G2F_ISR_TILE_6_F_LSB 6
`define GLC_STRM_G2F_ISR_TILE_6_F_MSB 6
`define GLC_STRM_G2F_ISR_TILE_7_F_LSB 7
`define GLC_STRM_G2F_ISR_TILE_7_F_MSB 7
`define GLC_STRM_G2F_ISR_TILE_8_F_LSB 8
`define GLC_STRM_G2F_ISR_TILE_8_F_MSB 8
`define GLC_STRM_G2F_ISR_TILE_9_F_LSB 9
`define GLC_STRM_G2F_ISR_TILE_9_F_MSB 9
`define GLC_STRM_G2F_ISR_TILE_10_F_LSB 10
`define GLC_STRM_G2F_ISR_TILE_10_F_MSB 10
`define GLC_STRM_G2F_ISR_TILE_11_F_LSB 11
`define GLC_STRM_G2F_ISR_TILE_11_F_MSB 11
`define GLC_STRM_G2F_ISR_TILE_12_F_LSB 12
`define GLC_STRM_G2F_ISR_TILE_12_F_MSB 12
`define GLC_STRM_G2F_ISR_TILE_13_F_LSB 13
`define GLC_STRM_G2F_ISR_TILE_13_F_MSB 13
`define GLC_STRM_G2F_ISR_TILE_14_F_LSB 14
`define GLC_STRM_G2F_ISR_TILE_14_F_MSB 14
`define GLC_STRM_G2F_ISR_TILE_15_F_LSB 15
`define GLC_STRM_G2F_ISR_TILE_15_F_MSB 15
`define GLC_PAR_CFG_G2F_ISR_R 'h38
`define GLC_PAR_CFG_G2F_ISR_R_LSB 0
`define GLC_PAR_CFG_G2F_ISR_R_MSB 15
`define GLC_PAR_CFG_G2F_ISR_TILE_0_F_LSB 0
`define GLC_PAR_CFG_G2F_ISR_TILE_0_F_MSB 0
`define GLC_PAR_CFG_G2F_ISR_TILE_1_F_LSB 1
`define GLC_PAR_CFG_G2F_ISR_TILE_1_F_MSB 1
`define GLC_PAR_CFG_G2F_ISR_TILE_2_F_LSB 2
`define GLC_PAR_CFG_G2F_ISR_TILE_2_F_MSB 2
`define GLC_PAR_CFG_G2F_ISR_TILE_3_F_LSB 3
`define GLC_PAR_CFG_G2F_ISR_TILE_3_F_MSB 3
`define GLC_PAR_CFG_G2F_ISR_TILE_4_F_LSB 4
`define GLC_PAR_CFG_G2F_ISR_TILE_4_F_MSB 4
`define GLC_PAR_CFG_G2F_ISR_TILE_5_F_LSB 5
`define GLC_PAR_CFG_G2F_ISR_TILE_5_F_MSB 5
`define GLC_PAR_CFG_G2F_ISR_TILE_6_F_LSB 6
`define GLC_PAR_CFG_G2F_ISR_TILE_6_F_MSB 6
`define GLC_PAR_CFG_G2F_ISR_TILE_7_F_LSB 7
`define GLC_PAR_CFG_G2F_ISR_TILE_7_F_MSB 7
`define GLC_PAR_CFG_G2F_ISR_TILE_8_F_LSB 8
`define GLC_PAR_CFG_G2F_ISR_TILE_8_F_MSB 8
`define GLC_PAR_CFG_G2F_ISR_TILE_9_F_LSB 9
`define GLC_PAR_CFG_G2F_ISR_TILE_9_F_MSB 9
`define GLC_PAR_CFG_G2F_ISR_TILE_10_F_LSB 10
`define GLC_PAR_CFG_G2F_ISR_TILE_10_F_MSB 10
`define GLC_PAR_CFG_G2F_ISR_TILE_11_F_LSB 11
`define GLC_PAR_CFG_G2F_ISR_TILE_11_F_MSB 11
`define GLC_PAR_CFG_G2F_ISR_TILE_12_F_LSB 12
`define GLC_PAR_CFG_G2F_ISR_TILE_12_F_MSB 12
`define GLC_PAR_CFG_G2F_ISR_TILE_13_F_LSB 13
`define GLC_PAR_CFG_G2F_ISR_TILE_13_F_MSB 13
`define GLC_PAR_CFG_G2F_ISR_TILE_14_F_LSB 14
`define GLC_PAR_CFG_G2F_ISR_TILE_14_F_MSB 14
`define GLC_PAR_CFG_G2F_ISR_TILE_15_F_LSB 15
`define GLC_PAR_CFG_G2F_ISR_TILE_15_F_MSB 15
`define GLC_GLOBAL_ISR_R 'h3c
`define GLC_GLOBAL_ISR_R_LSB 0
`define GLC_GLOBAL_ISR_R_MSB 2
`define GLC_GLOBAL_ISR_STRM_F2G_F_LSB 0
`define GLC_GLOBAL_ISR_STRM_F2G_F_MSB 0
`define GLC_GLOBAL_ISR_STRM_G2F_F_LSB 1
`define GLC_GLOBAL_ISR_STRM_G2F_F_MSB 1
`define GLC_GLOBAL_ISR_PAR_CFG_G2F_F_LSB 2
`define GLC_GLOBAL_ISR_PAR_CFG_G2F_F_MSB 2
`define GLC_CGRA_CONFIG_ADDR_R 'h40
`define GLC_CGRA_CONFIG_ADDR_R_LSB 0
`define GLC_CGRA_CONFIG_ADDR_R_MSB 31
`define GLC_CGRA_CONFIG_ADDR_ADDR_F_LSB 0
`define GLC_CGRA_CONFIG_ADDR_ADDR_F_MSB 31
`define GLC_CGRA_CONFIG_WR_DATA_R 'h44
`define GLC_CGRA_CONFIG_WR_DATA_R_LSB 0
`define GLC_CGRA_CONFIG_WR_DATA_R_MSB 31
`define GLC_CGRA_CONFIG_WR_DATA_DATA_F_LSB 0
`define GLC_CGRA_CONFIG_WR_DATA_DATA_F_MSB 31
`define GLC_CGRA_CONFIG_WRITE_R 'h48
`define GLC_CGRA_CONFIG_WRITE_R_LSB 0
`define GLC_CGRA_CONFIG_WRITE_R_MSB 31
`define GLC_CGRA_CONFIG_WRITE_CNT_F_LSB 0
`define GLC_CGRA_CONFIG_WRITE_CNT_F_MSB 31
`define GLC_CGRA_CONFIG_READ_R 'h4c
`define GLC_CGRA_CONFIG_READ_R_LSB 0
`define GLC_CGRA_CONFIG_READ_R_MSB 31
`define GLC_CGRA_CONFIG_READ_CNT_F_LSB 0
`define GLC_CGRA_CONFIG_READ_CNT_F_MSB 31
`define GLC_CGRA_CONFIG_RD_DATA_R 'h50
`define GLC_CGRA_CONFIG_RD_DATA_R_LSB 0
`define GLC_CGRA_CONFIG_RD_DATA_R_MSB 31
`define GLC_CGRA_CONFIG_RD_DATA_DATA_F_LSB 0
`define GLC_CGRA_CONFIG_RD_DATA_DATA_F_MSB 31
`define GLC_GLB_FLUSH_CROSSBAR_R 'h54
`define GLC_GLB_FLUSH_CROSSBAR_R_LSB 0
`define GLC_GLB_FLUSH_CROSSBAR_R_MSB 31
`define GLC_GLB_FLUSH_CROSSBAR_SEL_F_LSB 0
`define GLC_GLB_FLUSH_CROSSBAR_SEL_F_MSB 31
