`ifndef GARNET_PARAM
`define GARNET_PARAM

package header;

localparam int NUM_PRR = 8;
localparam int NUM_PRR_WIDTH = $clog2(NUM_PRR);

endpackage
`endif
