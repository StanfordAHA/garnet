module AN2D0BWP16P90 ( 
input logic  A, 
input logic  B, 
output logic  Z); 
assign Z = (A & B); 
endmodule  
