`define GLB_CFG_TILE_CTRL                   'h00
`define GLB_CFG_LATENCY                     'h04
`define GLB_CFG_ST_DMA_HEADER_0_VALIDATE    'h08
`define GLB_CFG_ST_DMA_HEADER_0_START_ADDR  'h0C
`define GLB_CFG_ST_DMA_HEADER_0_NUM_WORDS   'h10
`define GLB_CFG_ST_DMA_HEADER_1_VALIDATE    'h14
`define GLB_CFG_ST_DMA_HEADER_1_START_ADDR  'h18
`define GLB_CFG_ST_DMA_HEADER_1_NUM_WORDS   'h1C
`define GLB_CFG_ST_DMA_HEADER_2_VALIDATE    'h20
`define GLB_CFG_ST_DMA_HEADER_2_START_ADDR  'h24
`define GLB_CFG_ST_DMA_HEADER_2_NUM_WORDS   'h28
`define GLB_CFG_ST_DMA_HEADER_3_VALIDATE    'h2C
`define GLB_CFG_ST_DMA_HEADER_3_START_ADDR  'h30
`define GLB_CFG_ST_DMA_HEADER_3_NUM_WORDS   'h34
`define GLB_CFG_LD_DMA_HEADER_0_VALIDATE    'h38
`define GLB_CFG_LD_DMA_HEADER_0_START_ADDR  'h3C
`define GLB_CFG_LD_DMA_HEADER_0_ACTIVE_CTRL 'h40
`define GLB_CFG_LD_DMA_HEADER_0_ITER_CTRL_0 'h44
`define GLB_CFG_LD_DMA_HEADER_0_ITER_CTRL_1 'h48
`define GLB_CFG_LD_DMA_HEADER_0_ITER_CTRL_2 'h4C
`define GLB_CFG_LD_DMA_HEADER_0_ITER_CTRL_3 'h50
`define GLB_CFG_LD_DMA_HEADER_1_VALIDATE    'h54
`define GLB_CFG_LD_DMA_HEADER_1_START_ADDR  'h58
`define GLB_CFG_LD_DMA_HEADER_1_ACTIVE_CTRL 'h5C
`define GLB_CFG_LD_DMA_HEADER_1_ITER_CTRL_0 'h60
`define GLB_CFG_LD_DMA_HEADER_1_ITER_CTRL_1 'h64
`define GLB_CFG_LD_DMA_HEADER_1_ITER_CTRL_2 'h68
`define GLB_CFG_LD_DMA_HEADER_1_ITER_CTRL_3 'h6C
`define GLB_CFG_LD_DMA_HEADER_2_VALIDATE    'h70
`define GLB_CFG_LD_DMA_HEADER_2_START_ADDR  'h74
`define GLB_CFG_LD_DMA_HEADER_2_ACTIVE_CTRL 'h78
`define GLB_CFG_LD_DMA_HEADER_2_ITER_CTRL_0 'h7C
`define GLB_CFG_LD_DMA_HEADER_2_ITER_CTRL_1 'h80
`define GLB_CFG_LD_DMA_HEADER_2_ITER_CTRL_2 'h84
`define GLB_CFG_LD_DMA_HEADER_2_ITER_CTRL_3 'h88
`define GLB_CFG_LD_DMA_HEADER_3_VALIDATE    'h8C
`define GLB_CFG_LD_DMA_HEADER_3_START_ADDR  'h90
`define GLB_CFG_LD_DMA_HEADER_3_ACTIVE_CTRL 'h94
`define GLB_CFG_LD_DMA_HEADER_3_ITER_CTRL_0 'h98
`define GLB_CFG_LD_DMA_HEADER_3_ITER_CTRL_1 'h9C
`define GLB_CFG_LD_DMA_HEADER_3_ITER_CTRL_2 'hA0
`define GLB_CFG_LD_DMA_HEADER_3_ITER_CTRL_3 'hA4
`define GLB_CFG_PC_DMA_HEADER_0_START_ADDR  'hA8
`define GLB_CFG_PC_DMA_HEADER_0_NUM_CFG     'hAC
