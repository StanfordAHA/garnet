`ifndef GLOBAL_BUFFER_PARAM
`define GLOBAL_BUFFER_PARAM
package global_buffer_param;
localparam int NUM_PRR = 4;
localparam int NUM_CGRA_COLS = 8;
localparam int NUM_GLB_TILES = 4;
localparam int NUM_COLS_PER_GROUP = 4;
localparam int BANKS_PER_TILE = 2;
localparam int BANK_ADDR_WIDTH = 16;
localparam int BANK_DATA_WIDTH = 64;
localparam int CGRA_DATA_WIDTH = 16;
localparam int AXI_DATA_WIDTH = 32;
localparam int CGRA_AXI_ADDR_WIDTH = 13;
localparam int CGRA_AXI_DATA_WIDTH = 32;
localparam int CGRA_CFG_ADDR_WIDTH = 32;
localparam int CGRA_CFG_DATA_WIDTH = 32;
localparam int LOAD_DMA_FIFO_DEPTH = 16;
localparam int STORE_DMA_FIFO_DEPTH = 4;
localparam int MAX_NUM_CHAIN = 8;
localparam int ST_DMA_VALID_MODE_VALID = 0;
localparam int ST_DMA_VALID_MODE_READY_VALID = 1;
localparam int ST_DMA_VALID_MODE_STATIC = 2;
localparam int LD_DMA_VALID_MODE_STATIC = 0;
localparam int LD_DMA_VALID_MODE_VALID = 1;
localparam int LD_DMA_VALID_MODE_READY_VALID = 2;
localparam int LD_DMA_FLUSH_MODE_EXTERNAL = 0;
localparam int LD_DMA_FLUSH_MODE_INTERNAL = 1;
localparam int SRAM_MACRO_WORD_SIZE = 64;
localparam int SRAM_MACRO_MUX_SIZE = 8;
localparam int SRAM_MACRO_NUM_SUBARRAYS = 2;
localparam int NUM_PRR_WIDTH = 2;
localparam int TILE_SEL_ADDR_WIDTH = 2;
localparam int CGRA_PER_GLB = 2;
localparam int BANK_SEL_ADDR_WIDTH = 1;
localparam int BANK_STRB_WIDTH = 8;
localparam int BANK_BYTE_OFFSET = 3;
localparam int GLB_ADDR_WIDTH = 19;
localparam int CGRA_BYTE_OFFSET = 1;
localparam int AXI_ADDR_WIDTH = 12;
localparam int AXI_ADDR_REG_WIDTH = 8;
localparam int AXI_STRB_WIDTH = 4;
localparam int AXI_BYTE_OFFSET = 2;
localparam int MAX_NUM_CFG_WIDTH = 16;
localparam int NUM_GROUPS = 2;
localparam int QUEUE_DEPTH = 1;
localparam int LOAD_DMA_LOOP_LEVEL = 8;
localparam int STORE_DMA_LOOP_LEVEL = 7;
localparam int LOOP_LEVEL = 8;
localparam int CHAIN_LATENCY_OVERHEAD = 3;
localparam int LATENCY_WIDTH = 6;
localparam int PCFG_LATENCY_WIDTH = 6;
localparam int SRAM_MACRO_READ_LATENCY = 1;
localparam int GLB_DMA2BANK_DELAY = 1;
localparam int GLB_SW2BANK_PIPELINE_DEPTH = 0;
localparam int GLB_BANK2SW_PIPELINE_DEPTH = 1;
localparam int GLB_BANK_MEMORY_PIPELINE_DEPTH = 0;
localparam int SRAM_GEN_PIPELINE_DEPTH = 0;
localparam int SRAM_GEN_OUTPUT_PIPELINE_DEPTH = 0;
localparam int GLS_PIPELINE_DEPTH = 0;
localparam int TILE2SRAM_WR_DELAY = 1;
localparam int TILE2SRAM_RD_DELAY = 3;
localparam int BANKMUX2SRAM_WR_DELAY = 0;
localparam int BANKMUX2SRAM_RD_DELAY = 2;
localparam int FLUSH_CROSSBAR_PIPELINE_DEPTH = 1;
localparam int RD_CLK_EN_MARGIN = 3;
localparam int WR_CLK_EN_MARGIN = 3;
localparam int PROC_CLK_EN_MARGIN = 4;
localparam int IS_SRAM_STUB = 0;
localparam int CONFIG_PORT_PIPELINE_DEPTH = 1;
localparam int CYCLE_COUNT_WIDTH = 16;
localparam int INTERRUPT_CNT = 5;
endpackage
`endif
