`ifndef MATRIX_UNIT_PARAM
`define MATRIX_UNIT_PARAM
package matrix_unit_param;
localparam int MU_DATAWIDTH = 16;
localparam int OC_0 = 32;
endpackage
`endif
