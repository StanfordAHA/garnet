module global_buffer #(
    parameter integer BANK_DATA_WIDTH = 64,
    parameter integer CGRA_DATA_WIDTH = 16,
    parameter integer CFG_ADDR_WIDTH = 32,
    parameter integer CFG_DATA_WIDTH = 32,
    parameter integer GLB_CFG_ADDR_WIDTH = 12,
    parameter integer GLB_CFG_TILE_WIDTH = 2,
    parameter integer GLB_CFG_FEATURE_WIDTH = 4,
    parameter integer GLB_CFG_REG_WIDTH = 4,
    parameter integer BANK_ADDR_WIDTH = 17,
    parameter integer GLB_ADDR_WIDTH = 32
)
(
    input                                   clk,
    input                                   reset,

    input        [BANK_DATA_WIDTH/8-1:0]    host_wr_strb,
    input        [GLB_ADDR_WIDTH-1:0]       host_wr_addr,
    input        [BANK_DATA_WIDTH-1:0]      host_wr_data,

    input                                   host_rd_en,
    input        [GLB_ADDR_WIDTH-1:0]       host_rd_addr,
    output logic [BANK_DATA_WIDTH-1:0]      host_rd_data,

    input                                   cgra_to_io_wr_en [7:0],
    input                                   cgra_to_io_rd_en [7:0],
    output logic                            io_to_cgra_rd_data_valid [7:0],
    input        [CGRA_DATA_WIDTH-1:0]      cgra_to_io_wr_data [7:0],
    output logic [CGRA_DATA_WIDTH-1:0]      io_to_cgra_rd_data [7:0],
    input        [CGRA_DATA_WIDTH-1:0]      cgra_to_io_addr_high [7:0],
    input        [CGRA_DATA_WIDTH-1:0]      cgra_to_io_addr_low [7:0],

    input                                   glc_to_cgra_cfg_wr,
    input                                   glc_to_cgra_cfg_rd,
    input        [CFG_ADDR_WIDTH-1:0]       glc_to_cgra_cfg_addr,
    input        [CFG_DATA_WIDTH-1:0]       glc_to_cgra_cfg_data,

    output logic                            glb_to_cgra_cfg_wr [7:0],
    output logic                            glb_to_cgra_cfg_rd [7:0],
    output logic [CFG_ADDR_WIDTH-1:0]       glb_to_cgra_cfg_addr [7:0],
    output logic [CFG_DATA_WIDTH-1:0]       glb_to_cgra_cfg_data [7:0],

    input                                   glc_to_io_stall,
    input                                   cgra_start_pulse,
    output logic                            cgra_done_pulse,
    input                                   config_start_pulse,
    output logic                            config_done_pulse,

    input                                   glb_config_wr,
    input                                   glb_config_rd,
    input        [GLB_CFG_ADDR_WIDTH-1:0]   glb_config_addr,
    input        [CFG_DATA_WIDTH-1:0]       glb_config_wr_data,
    output logic [CFG_DATA_WIDTH-1:0]       glb_config_rd_data,

    input                                   glb_sram_config_wr,
    input                                   glb_sram_config_rd,
    input        [CFG_ADDR_WIDTH-1:0]       glb_sram_config_addr,
    input        [CFG_DATA_WIDTH-1:0]       glb_sram_config_wr_data,
    output logic [CFG_DATA_WIDTH-1:0]       glb_sram_config_rd_data
);
logic host_wr_en;
assign host_wr_en = |host_wr_strb;

    GlobalBuffer_32_8_8 glb_inst (
        .cgra_done_pulse(cgra_done_pulse),
        .cgra_start_pulse(cgra_start_pulse),
        .cgra_to_io_addr_high_0(cgra_to_io_addr_high[0]),
        .cgra_to_io_addr_high_1(cgra_to_io_addr_high[1]),
        .cgra_to_io_addr_high_2(cgra_to_io_addr_high[2]),
        .cgra_to_io_addr_high_3(cgra_to_io_addr_high[3]),
        .cgra_to_io_addr_high_4(cgra_to_io_addr_high[4]),
        .cgra_to_io_addr_high_5(cgra_to_io_addr_high[5]),
        .cgra_to_io_addr_high_6(cgra_to_io_addr_high[6]),
        .cgra_to_io_addr_high_7(cgra_to_io_addr_high[7]),
        .cgra_to_io_addr_low_0(cgra_to_io_addr_low[0]),
        .cgra_to_io_addr_low_1(cgra_to_io_addr_low[1]),
        .cgra_to_io_addr_low_2(cgra_to_io_addr_low[2]),
        .cgra_to_io_addr_low_3(cgra_to_io_addr_low[3]),
        .cgra_to_io_addr_low_4(cgra_to_io_addr_low[4]),
        .cgra_to_io_addr_low_5(cgra_to_io_addr_low[5]),
        .cgra_to_io_addr_low_6(cgra_to_io_addr_low[6]),
        .cgra_to_io_addr_low_7(cgra_to_io_addr_low[7]),
        .cgra_to_io_rd_en({cgra_to_io_rd_en[7],cgra_to_io_rd_en[6],  cgra_to_io_rd_en[5], cgra_to_io_rd_en[4], cgra_to_io_rd_en[3], cgra_to_io_rd_en[2], cgra_to_io_rd_en[1], cgra_to_io_rd_en[0]}),
        .cgra_to_io_wr_data_0(cgra_to_io_wr_data[0]),
        .cgra_to_io_wr_data_1(cgra_to_io_wr_data[1]),
        .cgra_to_io_wr_data_2(cgra_to_io_wr_data[2]),
        .cgra_to_io_wr_data_3(cgra_to_io_wr_data[3]),
        .cgra_to_io_wr_data_4(cgra_to_io_wr_data[4]),
        .cgra_to_io_wr_data_5(cgra_to_io_wr_data[5]),
        .cgra_to_io_wr_data_6(cgra_to_io_wr_data[6]),
        .cgra_to_io_wr_data_7(cgra_to_io_wr_data[7]),
        .cgra_to_io_wr_en({cgra_to_io_wr_en[7],cgra_to_io_wr_en[6],  cgra_to_io_wr_en[5], cgra_to_io_wr_en[4], cgra_to_io_wr_en[3], cgra_to_io_wr_en[2], cgra_to_io_wr_en[1], cgra_to_io_wr_en[0]}),
        .clk(clk),
        .config_done_pulse(config_done_pulse),
        .config_start_pulse(config_start_pulse),
        .glb_config_addr(glb_config_addr),
        .glb_config_rd(glb_config_rd),
        .glb_config_rd_data(glb_config_rd_data),
        .glb_config_wr(glb_config_wr),
        .glb_config_wr_data(glb_config_wr_data),
        .glb_sram_config_addr(glb_sram_config_addr),
        .glb_sram_config_rd(glb_sram_config_rd),
        .glb_sram_config_rd_data(glb_sram_config_rd_data),
        .glb_sram_config_wr(glb_sram_config_wr),
        .glb_sram_config_wr_data(glb_sram_config_wr_data),
        .glb_to_cgra_cfg_data_0(glb_to_cgra_cfg_data[0]),
        .glb_to_cgra_cfg_data_1(glb_to_cgra_cfg_data[1]),
        .glb_to_cgra_cfg_data_2(glb_to_cgra_cfg_data[2]),
        .glb_to_cgra_cfg_data_3(glb_to_cgra_cfg_data[3]),
        .glb_to_cgra_cfg_data_4(glb_to_cgra_cfg_data[4]),
        .glb_to_cgra_cfg_data_5(glb_to_cgra_cfg_data[5]),
        .glb_to_cgra_cfg_data_6(glb_to_cgra_cfg_data[6]),
        .glb_to_cgra_cfg_data_7(glb_to_cgra_cfg_data[7]),
        .glb_to_cgra_cfg_addr_0(glb_to_cgra_cfg_addr[0]),
        .glb_to_cgra_cfg_addr_1(glb_to_cgra_cfg_addr[1]),
        .glb_to_cgra_cfg_addr_2(glb_to_cgra_cfg_addr[2]),
        .glb_to_cgra_cfg_addr_3(glb_to_cgra_cfg_addr[3]),
        .glb_to_cgra_cfg_addr_4(glb_to_cgra_cfg_addr[4]),
        .glb_to_cgra_cfg_addr_5(glb_to_cgra_cfg_addr[5]),
        .glb_to_cgra_cfg_addr_6(glb_to_cgra_cfg_addr[6]),
        .glb_to_cgra_cfg_addr_7(glb_to_cgra_cfg_addr[7]),
        .glb_to_cgra_cfg_wr({glb_to_cgra_cfg_wr[7],glb_to_cgra_cfg_wr[6],  glb_to_cgra_cfg_wr[5], glb_to_cgra_cfg_wr[4], glb_to_cgra_cfg_wr[3], glb_to_cgra_cfg_wr[2], glb_to_cgra_cfg_wr[1], glb_to_cgra_cfg_wr[0]}),
        .glb_to_cgra_cfg_rd({glb_to_cgra_cfg_rd[7],glb_to_cgra_cfg_rd[6],  glb_to_cgra_cfg_rd[5], glb_to_cgra_cfg_rd[4], glb_to_cgra_cfg_rd[3], glb_to_cgra_cfg_rd[2], glb_to_cgra_cfg_rd[1], glb_to_cgra_cfg_rd[0]}),

        .glc_to_cgra_cfg_addr(glc_to_cgra_cfg_addr),
        .glc_to_cgra_cfg_data(glc_to_cgra_cfg_data),
        .glc_to_cgra_cfg_rd(glc_to_cgra_cfg_rd),
        .glc_to_cgra_cfg_wr(glc_to_cgra_cfg_wr),
        .host_rd_addr(host_rd_addr),
        .host_rd_data(host_rd_data),
        .host_rd_en(host_rd_en),
        .host_wr_addr(host_wr_addr),
        .host_wr_data(host_wr_data),
        .host_wr_en(host_wr_en),
        .host_wr_strb(host_wr_strb),
        .io_to_cgra_rd_data_0(io_to_cgra_rd_data[0]),
        .io_to_cgra_rd_data_1(io_to_cgra_rd_data[1]),
        .io_to_cgra_rd_data_2(io_to_cgra_rd_data[2]),
        .io_to_cgra_rd_data_3(io_to_cgra_rd_data[3]),
        .io_to_cgra_rd_data_4(io_to_cgra_rd_data[4]),
        .io_to_cgra_rd_data_5(io_to_cgra_rd_data[5]),
        .io_to_cgra_rd_data_6(io_to_cgra_rd_data[6]),
        .io_to_cgra_rd_data_7(io_to_cgra_rd_data[7]),
        .io_to_cgra_rd_data_valid({io_to_cgra_rd_data_valid[7],io_to_cgra_rd_data_valid[6],  io_to_cgra_rd_data_valid[5], io_to_cgra_rd_data_valid[4], io_to_cgra_rd_data_valid[3], io_to_cgra_rd_data_valid[2], io_to_cgra_rd_data_valid[1], io_to_cgra_rd_data_valid[0]}),
        .reset(reset),
        .stall(glc_to_io_stall)
    );

endmodule
