module pe_core
  (
   input [15:0]  data0,
   input [15:0]  data1,
   input [0:0]   bit0,
   input [0:0]   bit1,
   input [0:0]   bit2,
   output [15:0] res,
   output [0:0]  res_p
   );

endmodule
