module sink_64 (
    input logic[63:0] sink_in
); 
endmodule
