module SC7P5T_AN2X0P5_SSC14R ( 
input logic  A, 
input logic  B, 
output logic  Z); 
assign Z = (A & B); 
endmodule  
