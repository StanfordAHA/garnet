`define GLB_DATA_NETWORK_CTRL_R 'h0
`define GLB_DATA_NETWORK_CTRL_R_LSB 0
`define GLB_DATA_NETWORK_CTRL_R_MSB 0
`define GLB_DATA_NETWORK_CTRL_CONNECTED_F_LSB 0
`define GLB_DATA_NETWORK_CTRL_CONNECTED_F_MSB 0
`define GLB_DATA_NETWORK_LATENCY_R 'h4
`define GLB_DATA_NETWORK_LATENCY_R_LSB 0
`define GLB_DATA_NETWORK_LATENCY_R_MSB 5
`define GLB_DATA_NETWORK_LATENCY_VALUE_F_LSB 0
`define GLB_DATA_NETWORK_LATENCY_VALUE_F_MSB 5
`define GLB_PCFG_NETWORK_CTRL_R 'h8
`define GLB_PCFG_NETWORK_CTRL_R_LSB 0
`define GLB_PCFG_NETWORK_CTRL_R_MSB 0
`define GLB_PCFG_NETWORK_CTRL_CONNECTED_F_LSB 0
`define GLB_PCFG_NETWORK_CTRL_CONNECTED_F_MSB 0
`define GLB_PCFG_NETWORK_LATENCY_R 'hc
`define GLB_PCFG_NETWORK_LATENCY_R_LSB 0
`define GLB_PCFG_NETWORK_LATENCY_R_MSB 5
`define GLB_PCFG_NETWORK_LATENCY_VALUE_F_LSB 0
`define GLB_PCFG_NETWORK_LATENCY_VALUE_F_MSB 5
`define GLB_ST_DMA_CTRL_R 'h10
`define GLB_ST_DMA_CTRL_R_LSB 0
`define GLB_ST_DMA_CTRL_R_MSB 6
`define GLB_ST_DMA_CTRL_MODE_F_LSB 0
`define GLB_ST_DMA_CTRL_MODE_F_MSB 1
`define GLB_ST_DMA_CTRL_VALID_MODE_F_LSB 2
`define GLB_ST_DMA_CTRL_VALID_MODE_F_MSB 3
`define GLB_ST_DMA_CTRL_DATA_MUX_F_LSB 4
`define GLB_ST_DMA_CTRL_DATA_MUX_F_MSB 5
`define GLB_ST_DMA_CTRL_NUM_REPEAT_F_LSB 6
`define GLB_ST_DMA_CTRL_NUM_REPEAT_F_MSB 6
`define GLB_ST_DMA_NUM_BLOCKS_R 'h14
`define GLB_ST_DMA_NUM_BLOCKS_R_LSB 0
`define GLB_ST_DMA_NUM_BLOCKS_R_MSB 31
`define GLB_ST_DMA_NUM_BLOCKS_VALUE_F_LSB 0
`define GLB_ST_DMA_NUM_BLOCKS_VALUE_F_MSB 31
`define GLB_ST_DMA_RV_SEG_MODE_R 'h18
`define GLB_ST_DMA_RV_SEG_MODE_R_LSB 0
`define GLB_ST_DMA_RV_SEG_MODE_R_MSB 0
`define GLB_ST_DMA_RV_SEG_MODE_VALUE_F_LSB 0
`define GLB_ST_DMA_RV_SEG_MODE_VALUE_F_MSB 0
`define GLB_ST_DMA_HEADER_0_DIM_R 'h1c
`define GLB_ST_DMA_HEADER_0_DIM_R_LSB 0
`define GLB_ST_DMA_HEADER_0_DIM_R_MSB 3
`define GLB_ST_DMA_HEADER_0_DIM_DIM_F_LSB 0
`define GLB_ST_DMA_HEADER_0_DIM_DIM_F_MSB 3
`define GLB_ST_DMA_HEADER_0_START_ADDR_R 'h20
`define GLB_ST_DMA_HEADER_0_START_ADDR_R_LSB 0
`define GLB_ST_DMA_HEADER_0_START_ADDR_R_MSB 18
`define GLB_ST_DMA_HEADER_0_START_ADDR_START_ADDR_F_LSB 0
`define GLB_ST_DMA_HEADER_0_START_ADDR_START_ADDR_F_MSB 18
`define GLB_ST_DMA_HEADER_0_CYCLE_START_ADDR_R 'h24
`define GLB_ST_DMA_HEADER_0_CYCLE_START_ADDR_R_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_START_ADDR_R_MSB 15
`define GLB_ST_DMA_HEADER_0_CYCLE_START_ADDR_CYCLE_START_ADDR_F_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_START_ADDR_CYCLE_START_ADDR_F_MSB 15
`define GLB_ST_DMA_HEADER_0_RANGE_0_R 'h28
`define GLB_ST_DMA_HEADER_0_RANGE_0_R_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_0_R_MSB 31
`define GLB_ST_DMA_HEADER_0_RANGE_0_RANGE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_0_RANGE_F_MSB 31
`define GLB_ST_DMA_HEADER_0_STRIDE_0_R 'h2c
`define GLB_ST_DMA_HEADER_0_STRIDE_0_R_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_0_R_MSB 19
`define GLB_ST_DMA_HEADER_0_STRIDE_0_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_0_STRIDE_F_MSB 19
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_0_R 'h30
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_0_R_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_0_R_MSB 15
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_0_CYCLE_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_0_CYCLE_STRIDE_F_MSB 15
`define GLB_ST_DMA_HEADER_0_RANGE_1_R 'h34
`define GLB_ST_DMA_HEADER_0_RANGE_1_R_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_1_R_MSB 31
`define GLB_ST_DMA_HEADER_0_RANGE_1_RANGE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_1_RANGE_F_MSB 31
`define GLB_ST_DMA_HEADER_0_STRIDE_1_R 'h38
`define GLB_ST_DMA_HEADER_0_STRIDE_1_R_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_1_R_MSB 19
`define GLB_ST_DMA_HEADER_0_STRIDE_1_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_1_STRIDE_F_MSB 19
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_1_R 'h3c
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_1_R_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_1_R_MSB 15
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_1_CYCLE_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_1_CYCLE_STRIDE_F_MSB 15
`define GLB_ST_DMA_HEADER_0_RANGE_2_R 'h40
`define GLB_ST_DMA_HEADER_0_RANGE_2_R_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_2_R_MSB 31
`define GLB_ST_DMA_HEADER_0_RANGE_2_RANGE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_2_RANGE_F_MSB 31
`define GLB_ST_DMA_HEADER_0_STRIDE_2_R 'h44
`define GLB_ST_DMA_HEADER_0_STRIDE_2_R_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_2_R_MSB 19
`define GLB_ST_DMA_HEADER_0_STRIDE_2_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_2_STRIDE_F_MSB 19
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_2_R 'h48
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_2_R_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_2_R_MSB 15
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_2_CYCLE_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_2_CYCLE_STRIDE_F_MSB 15
`define GLB_ST_DMA_HEADER_0_RANGE_3_R 'h4c
`define GLB_ST_DMA_HEADER_0_RANGE_3_R_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_3_R_MSB 31
`define GLB_ST_DMA_HEADER_0_RANGE_3_RANGE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_3_RANGE_F_MSB 31
`define GLB_ST_DMA_HEADER_0_STRIDE_3_R 'h50
`define GLB_ST_DMA_HEADER_0_STRIDE_3_R_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_3_R_MSB 19
`define GLB_ST_DMA_HEADER_0_STRIDE_3_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_3_STRIDE_F_MSB 19
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_3_R 'h54
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_3_R_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_3_R_MSB 15
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_3_CYCLE_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_3_CYCLE_STRIDE_F_MSB 15
`define GLB_ST_DMA_HEADER_0_RANGE_4_R 'h58
`define GLB_ST_DMA_HEADER_0_RANGE_4_R_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_4_R_MSB 31
`define GLB_ST_DMA_HEADER_0_RANGE_4_RANGE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_4_RANGE_F_MSB 31
`define GLB_ST_DMA_HEADER_0_STRIDE_4_R 'h5c
`define GLB_ST_DMA_HEADER_0_STRIDE_4_R_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_4_R_MSB 19
`define GLB_ST_DMA_HEADER_0_STRIDE_4_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_4_STRIDE_F_MSB 19
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_4_R 'h60
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_4_R_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_4_R_MSB 15
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_4_CYCLE_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_4_CYCLE_STRIDE_F_MSB 15
`define GLB_ST_DMA_HEADER_0_RANGE_5_R 'h64
`define GLB_ST_DMA_HEADER_0_RANGE_5_R_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_5_R_MSB 31
`define GLB_ST_DMA_HEADER_0_RANGE_5_RANGE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_5_RANGE_F_MSB 31
`define GLB_ST_DMA_HEADER_0_STRIDE_5_R 'h68
`define GLB_ST_DMA_HEADER_0_STRIDE_5_R_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_5_R_MSB 19
`define GLB_ST_DMA_HEADER_0_STRIDE_5_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_5_STRIDE_F_MSB 19
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_5_R 'h6c
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_5_R_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_5_R_MSB 15
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_5_CYCLE_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_5_CYCLE_STRIDE_F_MSB 15
`define GLB_ST_DMA_HEADER_0_RANGE_6_R 'h70
`define GLB_ST_DMA_HEADER_0_RANGE_6_R_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_6_R_MSB 31
`define GLB_ST_DMA_HEADER_0_RANGE_6_RANGE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_RANGE_6_RANGE_F_MSB 31
`define GLB_ST_DMA_HEADER_0_STRIDE_6_R 'h74
`define GLB_ST_DMA_HEADER_0_STRIDE_6_R_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_6_R_MSB 19
`define GLB_ST_DMA_HEADER_0_STRIDE_6_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_STRIDE_6_STRIDE_F_MSB 19
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_6_R 'h78
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_6_R_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_6_R_MSB 15
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_6_CYCLE_STRIDE_F_LSB 0
`define GLB_ST_DMA_HEADER_0_CYCLE_STRIDE_6_CYCLE_STRIDE_F_MSB 15
`define GLB_LD_DMA_CTRL_R 'h7c
`define GLB_LD_DMA_CTRL_R_LSB 0
`define GLB_LD_DMA_CTRL_R_MSB 7
`define GLB_LD_DMA_CTRL_MODE_F_LSB 0
`define GLB_LD_DMA_CTRL_MODE_F_MSB 1
`define GLB_LD_DMA_CTRL_VALID_MODE_F_LSB 2
`define GLB_LD_DMA_CTRL_VALID_MODE_F_MSB 3
`define GLB_LD_DMA_CTRL_FLUSH_MODE_F_LSB 4
`define GLB_LD_DMA_CTRL_FLUSH_MODE_F_MSB 4
`define GLB_LD_DMA_CTRL_DATA_MUX_F_LSB 5
`define GLB_LD_DMA_CTRL_DATA_MUX_F_MSB 6
`define GLB_LD_DMA_CTRL_NUM_REPEAT_F_LSB 7
`define GLB_LD_DMA_CTRL_NUM_REPEAT_F_MSB 7
`define GLB_LD_DMA_HEADER_0_DIM_R 'h80
`define GLB_LD_DMA_HEADER_0_DIM_R_LSB 0
`define GLB_LD_DMA_HEADER_0_DIM_R_MSB 3
`define GLB_LD_DMA_HEADER_0_DIM_DIM_F_LSB 0
`define GLB_LD_DMA_HEADER_0_DIM_DIM_F_MSB 3
`define GLB_LD_DMA_HEADER_0_START_ADDR_R 'h84
`define GLB_LD_DMA_HEADER_0_START_ADDR_R_LSB 0
`define GLB_LD_DMA_HEADER_0_START_ADDR_R_MSB 18
`define GLB_LD_DMA_HEADER_0_START_ADDR_START_ADDR_F_LSB 0
`define GLB_LD_DMA_HEADER_0_START_ADDR_START_ADDR_F_MSB 18
`define GLB_LD_DMA_HEADER_0_CYCLE_START_ADDR_R 'h88
`define GLB_LD_DMA_HEADER_0_CYCLE_START_ADDR_R_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_START_ADDR_R_MSB 15
`define GLB_LD_DMA_HEADER_0_CYCLE_START_ADDR_CYCLE_START_ADDR_F_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_START_ADDR_CYCLE_START_ADDR_F_MSB 15
`define GLB_LD_DMA_HEADER_0_RANGE_0_R 'h8c
`define GLB_LD_DMA_HEADER_0_RANGE_0_R_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_0_R_MSB 31
`define GLB_LD_DMA_HEADER_0_RANGE_0_RANGE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_0_RANGE_F_MSB 31
`define GLB_LD_DMA_HEADER_0_STRIDE_0_R 'h90
`define GLB_LD_DMA_HEADER_0_STRIDE_0_R_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_0_R_MSB 19
`define GLB_LD_DMA_HEADER_0_STRIDE_0_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_0_STRIDE_F_MSB 19
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_0_R 'h94
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_0_R_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_0_R_MSB 15
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_0_CYCLE_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_0_CYCLE_STRIDE_F_MSB 15
`define GLB_LD_DMA_HEADER_0_RANGE_1_R 'h98
`define GLB_LD_DMA_HEADER_0_RANGE_1_R_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_1_R_MSB 31
`define GLB_LD_DMA_HEADER_0_RANGE_1_RANGE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_1_RANGE_F_MSB 31
`define GLB_LD_DMA_HEADER_0_STRIDE_1_R 'h9c
`define GLB_LD_DMA_HEADER_0_STRIDE_1_R_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_1_R_MSB 19
`define GLB_LD_DMA_HEADER_0_STRIDE_1_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_1_STRIDE_F_MSB 19
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_1_R 'ha0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_1_R_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_1_R_MSB 15
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_1_CYCLE_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_1_CYCLE_STRIDE_F_MSB 15
`define GLB_LD_DMA_HEADER_0_RANGE_2_R 'ha4
`define GLB_LD_DMA_HEADER_0_RANGE_2_R_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_2_R_MSB 31
`define GLB_LD_DMA_HEADER_0_RANGE_2_RANGE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_2_RANGE_F_MSB 31
`define GLB_LD_DMA_HEADER_0_STRIDE_2_R 'ha8
`define GLB_LD_DMA_HEADER_0_STRIDE_2_R_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_2_R_MSB 19
`define GLB_LD_DMA_HEADER_0_STRIDE_2_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_2_STRIDE_F_MSB 19
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_2_R 'hac
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_2_R_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_2_R_MSB 15
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_2_CYCLE_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_2_CYCLE_STRIDE_F_MSB 15
`define GLB_LD_DMA_HEADER_0_RANGE_3_R 'hb0
`define GLB_LD_DMA_HEADER_0_RANGE_3_R_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_3_R_MSB 31
`define GLB_LD_DMA_HEADER_0_RANGE_3_RANGE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_3_RANGE_F_MSB 31
`define GLB_LD_DMA_HEADER_0_STRIDE_3_R 'hb4
`define GLB_LD_DMA_HEADER_0_STRIDE_3_R_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_3_R_MSB 19
`define GLB_LD_DMA_HEADER_0_STRIDE_3_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_3_STRIDE_F_MSB 19
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_3_R 'hb8
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_3_R_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_3_R_MSB 15
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_3_CYCLE_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_3_CYCLE_STRIDE_F_MSB 15
`define GLB_LD_DMA_HEADER_0_RANGE_4_R 'hbc
`define GLB_LD_DMA_HEADER_0_RANGE_4_R_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_4_R_MSB 31
`define GLB_LD_DMA_HEADER_0_RANGE_4_RANGE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_4_RANGE_F_MSB 31
`define GLB_LD_DMA_HEADER_0_STRIDE_4_R 'hc0
`define GLB_LD_DMA_HEADER_0_STRIDE_4_R_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_4_R_MSB 19
`define GLB_LD_DMA_HEADER_0_STRIDE_4_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_4_STRIDE_F_MSB 19
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_4_R 'hc4
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_4_R_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_4_R_MSB 15
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_4_CYCLE_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_4_CYCLE_STRIDE_F_MSB 15
`define GLB_LD_DMA_HEADER_0_RANGE_5_R 'hc8
`define GLB_LD_DMA_HEADER_0_RANGE_5_R_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_5_R_MSB 31
`define GLB_LD_DMA_HEADER_0_RANGE_5_RANGE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_5_RANGE_F_MSB 31
`define GLB_LD_DMA_HEADER_0_STRIDE_5_R 'hcc
`define GLB_LD_DMA_HEADER_0_STRIDE_5_R_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_5_R_MSB 19
`define GLB_LD_DMA_HEADER_0_STRIDE_5_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_5_STRIDE_F_MSB 19
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_5_R 'hd0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_5_R_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_5_R_MSB 15
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_5_CYCLE_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_5_CYCLE_STRIDE_F_MSB 15
`define GLB_LD_DMA_HEADER_0_RANGE_6_R 'hd4
`define GLB_LD_DMA_HEADER_0_RANGE_6_R_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_6_R_MSB 31
`define GLB_LD_DMA_HEADER_0_RANGE_6_RANGE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_6_RANGE_F_MSB 31
`define GLB_LD_DMA_HEADER_0_STRIDE_6_R 'hd8
`define GLB_LD_DMA_HEADER_0_STRIDE_6_R_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_6_R_MSB 19
`define GLB_LD_DMA_HEADER_0_STRIDE_6_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_6_STRIDE_F_MSB 19
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_6_R 'hdc
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_6_R_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_6_R_MSB 15
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_6_CYCLE_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_6_CYCLE_STRIDE_F_MSB 15
`define GLB_LD_DMA_HEADER_0_RANGE_7_R 'he0
`define GLB_LD_DMA_HEADER_0_RANGE_7_R_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_7_R_MSB 31
`define GLB_LD_DMA_HEADER_0_RANGE_7_RANGE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_RANGE_7_RANGE_F_MSB 31
`define GLB_LD_DMA_HEADER_0_STRIDE_7_R 'he4
`define GLB_LD_DMA_HEADER_0_STRIDE_7_R_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_7_R_MSB 19
`define GLB_LD_DMA_HEADER_0_STRIDE_7_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_STRIDE_7_STRIDE_F_MSB 19
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_7_R 'he8
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_7_R_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_7_R_MSB 15
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_7_CYCLE_STRIDE_F_LSB 0
`define GLB_LD_DMA_HEADER_0_CYCLE_STRIDE_7_CYCLE_STRIDE_F_MSB 15
`define GLB_PCFG_DMA_CTRL_R 'hec
`define GLB_PCFG_DMA_CTRL_R_LSB 0
`define GLB_PCFG_DMA_CTRL_R_MSB 17
`define GLB_PCFG_DMA_CTRL_MODE_F_LSB 0
`define GLB_PCFG_DMA_CTRL_MODE_F_MSB 0
`define GLB_PCFG_DMA_CTRL_RELOCATION_VALUE_F_LSB 1
`define GLB_PCFG_DMA_CTRL_RELOCATION_VALUE_F_MSB 16
`define GLB_PCFG_DMA_CTRL_RELOCATION_IS_MSB_F_LSB 17
`define GLB_PCFG_DMA_CTRL_RELOCATION_IS_MSB_F_MSB 17
`define GLB_PCFG_DMA_HEADER_START_ADDR_R 'hf0
`define GLB_PCFG_DMA_HEADER_START_ADDR_R_LSB 0
`define GLB_PCFG_DMA_HEADER_START_ADDR_R_MSB 18
`define GLB_PCFG_DMA_HEADER_START_ADDR_START_ADDR_F_LSB 0
`define GLB_PCFG_DMA_HEADER_START_ADDR_START_ADDR_F_MSB 18
`define GLB_PCFG_DMA_HEADER_NUM_CFG_R 'hf4
`define GLB_PCFG_DMA_HEADER_NUM_CFG_R_LSB 0
`define GLB_PCFG_DMA_HEADER_NUM_CFG_R_MSB 15
`define GLB_PCFG_DMA_HEADER_NUM_CFG_NUM_CFG_F_LSB 0
`define GLB_PCFG_DMA_HEADER_NUM_CFG_NUM_CFG_F_MSB 15
`define GLB_PCFG_BROADCAST_MUX_R 'hf8
`define GLB_PCFG_BROADCAST_MUX_R_LSB 0
`define GLB_PCFG_BROADCAST_MUX_R_MSB 5
`define GLB_PCFG_BROADCAST_MUX_WEST_F_LSB 0
`define GLB_PCFG_BROADCAST_MUX_WEST_F_MSB 1
`define GLB_PCFG_BROADCAST_MUX_EAST_F_LSB 2
`define GLB_PCFG_BROADCAST_MUX_EAST_F_MSB 3
`define GLB_PCFG_BROADCAST_MUX_SOUTH_F_LSB 4
`define GLB_PCFG_BROADCAST_MUX_SOUTH_F_MSB 5
