module dummy();
endmodule
