module AN2D0BWP16P90 ( 
input logic  A1, 
input logic  A2, 
output logic  Z); 
assign Z = (A1 & A2); 
endmodule  
