`define GLC_TEST 'h0
`define GLC_GLOBAL_RESET 'h4
`define GLC_SOFT_RESET 'h8
`define GLC_STALL 'hc
`define GLC_STREAM_START_PULSE 'h10
`define GLC_PC_START_PULSE 'h14
`define GLC_STRM_F2G_IER 'h18
`define GLC_STRM_G2F_IER 'h1c
`define GLC_PAR_CFG_G2F_IER 'h20
`define GLC_GLOBAL_IER 'h24
`define GLC_STRM_F2G_ISR 'h28
`define GLC_STRM_G2F_ISR 'h2c
`define GLC_PAR_CFG_G2F_ISR 'h30
`define GLC_GLOBAL_ISR 'h34
`define GLC_CGRA_CONFIG 'h38
`define GLC_CGRA_CONFIG_ADDR 'h38
`define GLC_CGRA_CONFIG_WR_DATA 'h3c
`define GLC_CGRA_CONFIG_WRITE 'h40
`define GLC_CGRA_CONFIG_READ 'h44
`define GLC_CGRA_CONFIG_RD_DATA 'h48
