/*=============================================================================
** Module: io_address_generator.sv
** Description:
**              Address generator for I/O controller
** Author: Taeyoung Kong
** Change history: 04/10/2019 - Implement first version only with interface 
**                 05/10/2019 - INSTREAM, OUTSTREAM modes are implemented
**===========================================================================*/
import global_buffer_pkg::*;

module glb_fbrc_address_generator (
    input  logic                            clk,
    input  logic                            clk_en,
    input  logic                            reset,
    input  logic                            cgra_start_pulse,
    output logic                            cgra_done_pulse,

    input  logic [GLB_ADDR_WIDTH-1:0]       start_addr,
    input  logic [GLB_ADDR_WIDTH-1:0]       num_words,
    input  addr_gen_mode_t                  mode,
    input  logic [CONFIG_DATA_WIDTH-1:0]    done_delay,

    input  logic                            cgra_to_io_wr_en,
    input  logic                            cgra_to_io_rd_en,
    input  logic [CGRA_DATA_WIDTH-1:0]      cgra_to_io_wr_data,
    output logic [CGRA_DATA_WIDTH-1:0]      io_to_cgra_rd_data,
    output logic                            io_to_cgra_rd_data_valid,
    input  logic [CGRA_DATA_WIDTH-1:0]      cgra_to_io_addr_high,
    input  logic [CGRA_DATA_WIDTH-1:0]      cgra_to_io_addr_low,
    
    output logic                            io_to_bank_wr_en,
    output logic [BANK_DATA_WIDTH-1:0]      io_to_bank_wr_data,
    output logic [BANK_DATA_WIDTH-1:0]      io_to_bank_wr_data_bit_sel,
    output logic                            io_to_bank_rd_en,
    input  logic [BANK_DATA_WIDTH-1:0]      bank_to_io_rd_data,
    input  logic                            bank_to_io_rd_data_valid,
    output logic [GLB_ADDR_WIDTH-1:0]       io_to_bank_addr
);

//============================================================================//
// local parameter declaration
//============================================================================//
localparam integer DATA_SEL_WIDTH = $clog2(BANK_DATA_WIDTH/CGRA_DATA_WIDTH); //2
localparam integer CGRA_DATA_BYTE = ((CGRA_DATA_WIDTH + 8 - 1)/8); //2
localparam integer BANK_ADDR_OFFSET = $clog2(BANK_DATA_WIDTH/8); // 3

//============================================================================//
// register to latch data from bank
//============================================================================//
logic                       io_to_bank_rd_en_d1; 
logic                       io_to_bank_rd_en_d2; 
logic [BANK_DATA_WIDTH-1:0] bank_to_io_rd_data_reg;
logic                       bank_to_io_rd_data_valid_reg;
logic [BANK_DATA_WIDTH-1:0] int_bank_to_io_rd_data;
logic                       int_bank_to_io_rd_data_valid;

always_ff @(posedge clk) begin
    if (clk_en) begin
        io_to_bank_rd_en_d1 <= io_to_bank_rd_en;
        io_to_bank_rd_en_d2 <= io_to_bank_rd_en_d1;
        bank_to_io_rd_data_reg <= int_bank_to_io_rd_data;
        bank_to_io_rd_data_valid_reg <= int_bank_to_io_rd_data_valid;
    end
end
assign int_bank_to_io_rd_data = io_to_bank_rd_en_d2 ? bank_to_io_rd_data : bank_to_io_rd_data_reg;
assign int_bank_to_io_rd_data_valid = io_to_bank_rd_en_d2 ? bank_to_io_rd_data_valid : bank_to_io_rd_data_valid_reg;

//============================================================================//
// INSTREAM mode
//============================================================================//
enum logic[1:0] {IDLE_INSTREAM, READ_INSTREAM, DONE_INSTREAM} state_instream;

logic [GLB_ADDR_WIDTH-1:0]      int_addr_instream;

logic [GLB_ADDR_WIDTH-1:0]      num_words_cnt_instream;
logic [CONFIG_DATA_WIDTH-1:0]   done_cnt_instream;

logic [DATA_SEL_WIDTH-1:0]      data_sel_instream;
logic [DATA_SEL_WIDTH-1:0]      data_sel_instream_d1;
logic [DATA_SEL_WIDTH-1:0]      data_sel_instream_d2;

logic                           int_rd_data_valid_instream;
logic                           int_rd_data_valid_instream_d1;
logic                           int_rd_data_valid_instream_d2;

logic                           io_to_cgra_rd_data_valid_instream;
logic [CGRA_DATA_WIDTH-1:0]     io_to_cgra_rd_data_instream;

logic                           io_to_bank_rd_en_instream;
logic [GLB_ADDR_WIDTH-1:0]      io_to_bank_addr_instream;

logic                           cgra_done_pulse_instream;

// Need mux to select CGRA_DATA from BANK_DATA due to DATA_WIDTH difference
assign data_sel_instream = int_addr_instream[CGRA_DATA_BYTE-1 +: DATA_SEL_WIDTH];

// in INSTREAM mode, io_to_bank_addr is equal to
// int_addr_instream with ADDR_OFFSET bits set to 0
assign io_to_bank_addr_instream = {int_addr_instream[GLB_ADDR_WIDTH-1:BANK_ADDR_OFFSET], {BANK_ADDR_OFFSET{1'b0}}};

// FSM for INSTREAM mode
// address increases by CGRA_DATA_BYTE if num_words_cnt is greater than 1
// num_words_cnt decreases by 1 if it is non-zero
always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
        state_instream <= IDLE_INSTREAM;
        num_words_cnt_instream <= 0;
        done_cnt_instream <= 0;
        int_addr_instream <= 0;
        io_to_bank_rd_en_instream <= 0;
        cgra_done_pulse_instream <= 0;
    end
    else if (clk_en) begin
        if (mode == INSTREAM) begin
            if (cgra_start_pulse) begin
                if (num_words > 0) begin
                    state_instream <= READ_INSTREAM;
                    num_words_cnt_instream <= num_words;
                    done_cnt_instream <= done_delay;
                    int_addr_instream <= start_addr;
                    io_to_bank_rd_en_instream <= 1;
                    cgra_done_pulse_instream <= 0;
                end
                // corner case when num_words is set to 0 when cgra_start_pulse is high
                else begin
                    state_instream <= DONE_INSTREAM;
                    num_words_cnt_instream <= 0;
                    done_cnt_instream <= done_delay;
                    int_addr_instream <= start_addr;
                    io_to_bank_rd_en_instream <= 0;
                    cgra_done_pulse_instream <= 0;
                end
            end
            else begin
                case (state_instream)
                    IDLE_INSTREAM: begin
                        state_instream <= IDLE_INSTREAM;
                        num_words_cnt_instream <= 0;
                        done_cnt_instream <= 0;
                        int_addr_instream <= int_addr_instream;
                        io_to_bank_rd_en_instream <= 0;
                        cgra_done_pulse_instream <= 0;
                    end
                    READ_INSTREAM: begin
                        if (num_words_cnt_instream == 1) begin
                            state_instream <= DONE_INSTREAM;
                            num_words_cnt_instream <= 0;
                            done_cnt_instream <= done_cnt_instream;
                            int_addr_instream <= int_addr_instream;
                            io_to_bank_rd_en_instream <= 0;
                            cgra_done_pulse_instream <= 0;
                        end
                        else begin
                            state_instream <= READ_INSTREAM;
                            num_words_cnt_instream <= num_words_cnt_instream - 1;
                            done_cnt_instream <= done_cnt_instream;
                            int_addr_instream <= int_addr_instream + CGRA_DATA_BYTE;
                            // bank_rd_en goes high only when the last word is read
                            io_to_bank_rd_en_instream <= (data_sel_instream == {DATA_SEL_WIDTH{1'b1}});
                            cgra_done_pulse_instream <= 0;
                        end
                    end
                    DONE_INSTREAM: begin
                        if (done_cnt_instream == 0) begin
                            state_instream <= IDLE_INSTREAM;
                            num_words_cnt_instream <= 0;
                            done_cnt_instream <= 0;
                            int_addr_instream <= int_addr_instream;
                            io_to_bank_rd_en_instream <= 0;
                            cgra_done_pulse_instream <= 1;
                        end
                        else begin
                            state_instream <= DONE_INSTREAM;
                            num_words_cnt_instream <= 0;
                            done_cnt_instream <= done_cnt_instream - 1;
                            int_addr_instream <= int_addr_instream;
                            io_to_bank_rd_en_instream <= 0;
                            cgra_done_pulse_instream <= 0;
                        end
                    end
                    default: begin
                        state_instream <= IDLE_INSTREAM;
                        num_words_cnt_instream <= 0;
                        done_cnt_instream <= 0;
                        int_addr_instream <= int_addr_instream;
                        io_to_bank_rd_en_instream <= 0;
                        cgra_done_pulse_instream <= 0;
                    end
                endcase
            end
        end
        // Mode is not INSTREAM
        else begin
            state_instream <= IDLE_INSTREAM;
            num_words_cnt_instream <= 0;
            done_cnt_instream <= 0;
            int_addr_instream <= int_addr_instream;
            io_to_bank_rd_en_instream <= 0;
            cgra_done_pulse_instream <= 0;
        end
    end
end

// When num_words_cnt is non-zero, rd_data_valid is positive
// io_to_cgra_rd_data_valid goes high 2 cycles after num_cnt is greater than 0
// due to read latency
assign int_rd_data_valid_instream = (num_words_cnt_instream > 0);
always_ff @(posedge clk) begin
    if (clk_en) begin
        int_rd_data_valid_instream_d1 <= int_rd_data_valid_instream;
        int_rd_data_valid_instream_d2 <= int_rd_data_valid_instream_d1;
    end
end
assign io_to_cgra_rd_data_valid_instream = int_bank_to_io_rd_data_valid & int_rd_data_valid_instream_d2;

// Need mux to select CGRA_DATA from BANK_DATA due to DATA_WIDTH difference
always_ff @(posedge clk) begin
    if (clk_en) begin
        data_sel_instream_d1 <= data_sel_instream;
        data_sel_instream_d2 <= data_sel_instream_d1;
    end
end
assign io_to_cgra_rd_data_instream = int_bank_to_io_rd_data[data_sel_instream_d2 * CGRA_DATA_WIDTH +: CGRA_DATA_WIDTH];

//============================================================================//
// OUTSTREAM mode
//============================================================================//
enum logic[1:0] {IDLE_OUTSTREAM, WRITE_OUTSTREAM, DONE_OUTSTREAM} state_outstream;

logic [GLB_ADDR_WIDTH-1:0]      int_addr_outstream;

logic [GLB_ADDR_WIDTH-1:0]      num_words_cnt_outstream;
logic [CONFIG_DATA_WIDTH-1:0]   done_cnt_outstream;

logic                           io_to_bank_wr_en_outstream;
logic [BANK_DATA_WIDTH-1:0]     io_to_bank_wr_data_outstream;
logic [GLB_ADDR_WIDTH-1:0]      io_to_bank_addr_outstream;
logic [BANK_DATA_WIDTH-1:0]     io_to_bank_bit_sel_outstream;

logic                           cgra_to_io_wr_en_outstream;
logic [CGRA_DATA_WIDTH-1:0]     cgra_to_io_wr_data_outstream;

logic                           cgra_done_pulse_outstream;

logic [DATA_SEL_WIDTH-1:0]      data_sel_outstream;

// In OUTSTREAM mode, wr_en and wr_data comes from cgra
assign cgra_to_io_wr_en_outstream = cgra_to_io_wr_en;
assign cgra_to_io_wr_data_outstream = cgra_to_io_wr_data;
                                                 
// We need mux due to the difference BANK_DATA_WIDTH and CGRA_DATA_WIDTH
// It will be used to decide io_to_bank_bit_sel for partial write
assign data_sel_outstream = int_addr_outstream[CGRA_DATA_BYTE-1 +: DATA_SEL_WIDTH];

// FSM for OUTSTREAM mode
// address increases by CGRA_DATA_BYTE if num_words_cnt is greater than 1
// num_words_cnt decreases by 1 if it is non-zero
always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
        num_words_cnt_outstream <= 0;
        done_cnt_outstream <= 0;
        int_addr_outstream <= 0;
        state_outstream <= IDLE_OUTSTREAM;
        io_to_bank_wr_en_outstream <= 0;
        io_to_bank_wr_data_outstream <= 0;
        io_to_bank_addr_outstream <= 0;
        io_to_bank_bit_sel_outstream <= 0;
        cgra_done_pulse_outstream <= 0;
    end
    else if (clk_en) begin
        if (mode == OUTSTREAM) begin
            if (cgra_start_pulse) begin
                if (num_words > 0) begin
                    state_outstream <= WRITE_OUTSTREAM;
                    num_words_cnt_outstream <= num_words;
                    done_cnt_outstream <= done_delay;
                    int_addr_outstream <= start_addr;
                    io_to_bank_wr_en_outstream <= 0;
                    io_to_bank_wr_data_outstream <= 0;
                    io_to_bank_addr_outstream <= 0;
                    io_to_bank_bit_sel_outstream <= 0;
                    cgra_done_pulse_outstream <= 0;
                end
                else begin
                    state_outstream <= DONE_OUTSTREAM;
                    num_words_cnt_outstream <= 0;
                    done_cnt_outstream <= done_delay;
                    int_addr_outstream <= start_addr;
                    io_to_bank_wr_en_outstream <= 0;
                    io_to_bank_wr_data_outstream <= 0;
                    io_to_bank_addr_outstream <= 0;
                    io_to_bank_bit_sel_outstream <= 0;
                    cgra_done_pulse_outstream <= 0;
                end
            end
            else begin
                case (state_outstream)
                    IDLE_OUTSTREAM: begin
                        state_outstream <= IDLE_OUTSTREAM;
                        num_words_cnt_outstream <= 0;
                        done_cnt_outstream <= 0;
                        int_addr_outstream <= int_addr_outstream;
                        io_to_bank_wr_en_outstream <= 0;
                        io_to_bank_wr_data_outstream <= 0;
                        io_to_bank_addr_outstream <= 0;
                        io_to_bank_bit_sel_outstream <= 0;
                        cgra_done_pulse_outstream <= 0;
                    end
                    WRITE_OUTSTREAM: begin
                        if (cgra_to_io_wr_en_outstream) begin
                            if (num_words_cnt_outstream == 1) begin
                                state_outstream <= DONE_OUTSTREAM;
                                num_words_cnt_outstream <= 0;
                                done_cnt_outstream <= done_cnt_outstream;
                                int_addr_outstream <= int_addr_outstream;
                                io_to_bank_wr_en_outstream <= 1;
                                io_to_bank_wr_data_outstream[data_sel_outstream*CGRA_DATA_WIDTH +: CGRA_DATA_WIDTH] <= cgra_to_io_wr_data_outstream;
                                io_to_bank_bit_sel_outstream[data_sel_outstream*CGRA_DATA_WIDTH +: CGRA_DATA_WIDTH] <= {CGRA_DATA_WIDTH{1'b1}};
                                io_to_bank_addr_outstream <= {int_addr_outstream[GLB_ADDR_WIDTH-1:BANK_ADDR_OFFSET], {BANK_ADDR_OFFSET{1'b0}}};
                                cgra_done_pulse_outstream <= 0;
                            end
                            else if (data_sel_outstream == {DATA_SEL_WIDTH{1'b1}}) begin
                                state_outstream <= WRITE_OUTSTREAM;
                                num_words_cnt_outstream <= num_words_cnt_outstream - 1;
                                done_cnt_outstream <= done_cnt_outstream;
                                int_addr_outstream <= int_addr_outstream + CGRA_DATA_BYTE;
                                io_to_bank_wr_en_outstream <= 1;
                                io_to_bank_wr_data_outstream[data_sel_outstream*CGRA_DATA_WIDTH +: CGRA_DATA_WIDTH] <= cgra_to_io_wr_data_outstream;
                                io_to_bank_bit_sel_outstream[data_sel_outstream*CGRA_DATA_WIDTH +: CGRA_DATA_WIDTH] <= {CGRA_DATA_WIDTH{1'b1}};
                                io_to_bank_addr_outstream <= {int_addr_outstream[GLB_ADDR_WIDTH-1:BANK_ADDR_OFFSET], {BANK_ADDR_OFFSET{1'b0}}};
                                cgra_done_pulse_outstream <= 0;
                            end
                            else if (data_sel_outstream == {DATA_SEL_WIDTH{1'b0}}) begin
                                state_outstream <= WRITE_OUTSTREAM;
                                num_words_cnt_outstream <= num_words_cnt_outstream - 1;
                                done_cnt_outstream <= done_cnt_outstream;
                                int_addr_outstream <= int_addr_outstream + CGRA_DATA_BYTE;
                                io_to_bank_wr_en_outstream <= 0;
                                io_to_bank_wr_data_outstream[data_sel_outstream*CGRA_DATA_WIDTH +: CGRA_DATA_WIDTH] <= cgra_to_io_wr_data_outstream;
                                io_to_bank_bit_sel_outstream <= {{(BANK_DATA_WIDTH-CGRA_DATA_WIDTH){1'b0}}, {CGRA_DATA_WIDTH{1'b1}}};
                                io_to_bank_addr_outstream <= io_to_bank_addr_outstream;
                                cgra_done_pulse_outstream <= 0;
                            end
                            else begin
                                state_outstream <= WRITE_OUTSTREAM;
                                num_words_cnt_outstream <= num_words_cnt_outstream - 1;
                                done_cnt_outstream <= done_cnt_outstream;
                                int_addr_outstream <= int_addr_outstream + CGRA_DATA_BYTE;
                                io_to_bank_wr_en_outstream <= 0;
                                io_to_bank_wr_data_outstream[data_sel_outstream*CGRA_DATA_WIDTH +: CGRA_DATA_WIDTH] <= cgra_to_io_wr_data_outstream;
                                io_to_bank_bit_sel_outstream[data_sel_outstream*CGRA_DATA_WIDTH +: CGRA_DATA_WIDTH] <= {CGRA_DATA_WIDTH{1'b1}};
                                io_to_bank_addr_outstream <= io_to_bank_addr_outstream;
                                cgra_done_pulse_outstream <= 0;
                            end
                        end
                        else begin
                            state_outstream <= WRITE_OUTSTREAM;
                            num_words_cnt_outstream <= num_words_cnt_outstream;
                            done_cnt_outstream <= done_cnt_outstream;
                            int_addr_outstream <= int_addr_outstream;
                            io_to_bank_wr_en_outstream <= 0;
                            io_to_bank_wr_data_outstream <= io_to_bank_wr_data_outstream;
                            io_to_bank_bit_sel_outstream <= io_to_bank_bit_sel_outstream;
                            io_to_bank_addr_outstream <= io_to_bank_addr_outstream;
                            cgra_done_pulse_outstream <= 0;
                        end
                    end
                    DONE_OUTSTREAM: begin
                        if (done_cnt_outstream == 0) begin
                            state_outstream <= IDLE_OUTSTREAM;
                            num_words_cnt_outstream <= 0;
                            done_cnt_outstream <= 0;
                            int_addr_outstream <= int_addr_outstream;
                            io_to_bank_wr_en_outstream <= 0;
                            io_to_bank_wr_data_outstream <= io_to_bank_wr_data_outstream;
                            io_to_bank_bit_sel_outstream <= 0;
                            io_to_bank_addr_outstream <= io_to_bank_addr_outstream;
                            cgra_done_pulse_outstream <= 1;
                        end
                        else begin
                            state_outstream <= DONE_OUTSTREAM;
                            num_words_cnt_outstream <= 0;
                            done_cnt_outstream <= done_cnt_outstream - 1;
                            int_addr_outstream <= int_addr_outstream;
                            io_to_bank_wr_en_outstream <= 0;
                            io_to_bank_wr_data_outstream <= io_to_bank_wr_data_outstream;
                            io_to_bank_bit_sel_outstream <= 0;
                            io_to_bank_addr_outstream <= io_to_bank_addr_outstream;
                            cgra_done_pulse_outstream <= 0;
                        end
                    end
                    default: begin
                        state_outstream <= IDLE_OUTSTREAM;
                        num_words_cnt_outstream <= 0;
                        done_cnt_outstream <= done_cnt_outstream;
                        int_addr_outstream <= int_addr_outstream;
                        io_to_bank_wr_en_outstream <= 0;
                        io_to_bank_wr_data_outstream <= io_to_bank_wr_data_outstream;
                        io_to_bank_bit_sel_outstream <= 0;
                        io_to_bank_addr_outstream <= io_to_bank_addr_outstream;
                        cgra_done_pulse_outstream <= 0;
                    end
                endcase
            end
        end
        else begin
            state_outstream <= IDLE_OUTSTREAM;
            num_words_cnt_outstream <= 0;
            done_cnt_outstream <= 0;
            int_addr_outstream <= int_addr_outstream;
            io_to_bank_wr_en_outstream <= 0;
            io_to_bank_wr_data_outstream <= io_to_bank_wr_data_outstream;
            io_to_bank_bit_sel_outstream <= 0;
            io_to_bank_addr_outstream <= io_to_bank_addr_outstream;
            cgra_done_pulse_outstream <= 0;
        end
    end
end

//============================================================================//
// SRAM mode
// If num_words is set to n, it generates cgra_done_pulse when the sum of
// the number of cgra writes and reads becomes n.
// If both cgra_to_io_wr_en and cgra_to_io_rd_en are asserted at the same
// cycle (which is not desired scenario), cgra_to_io_wr_en has priority. 
//============================================================================//
enum logic[1:0] {IDLE_SRAM, RUN_SRAM, RUN_SRAM_LOOP, DONE_SRAM} state_sram;

logic [GLB_ADDR_WIDTH-1:0]      int_addr_sram;

logic [GLB_ADDR_WIDTH-1:0]      num_words_cnt_sram;
logic [CONFIG_DATA_WIDTH-1:0]   done_cnt_sram;

logic                           io_to_bank_wr_en_sram;
logic [BANK_DATA_WIDTH-1:0]     io_to_bank_wr_data_sram;
logic [GLB_ADDR_WIDTH-1:0]      io_to_bank_addr_sram;
logic [BANK_DATA_WIDTH-1:0]     io_to_bank_bit_sel_sram;
logic                           io_to_bank_rd_en_sram;
logic                           io_to_bank_rd_en_sram_d1;
logic                           io_to_bank_rd_en_sram_d2;

logic                           cgra_to_io_wr_en_sram;
logic                           cgra_to_io_rd_en_sram;
logic [CGRA_DATA_WIDTH-1:0]     cgra_to_io_wr_data_sram;
logic [CGRA_DATA_WIDTH-1:0]     io_to_cgra_rd_data_sram;
logic                           io_to_cgra_rd_data_valid_sram;

logic                           cgra_done_pulse_sram;

logic [DATA_SEL_WIDTH-1:0]      data_sel_sram;
logic [DATA_SEL_WIDTH-1:0]      data_sel_sram_d1;
logic [DATA_SEL_WIDTH-1:0]      data_sel_sram_d2;

// In SRAM mode, wr_en and wr_data comes from cgra
assign cgra_to_io_wr_en_sram = cgra_to_io_wr_en;
assign cgra_to_io_wr_data_sram = cgra_to_io_wr_data;
                                                 
// In SRAM mode, rd_en comes from cgra
assign cgra_to_io_rd_en_sram = cgra_to_io_rd_en;

// FSM for SRAM mode
// if num_words is set to 0, it does not generate cgra_done_pulse
always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
        state_sram <= IDLE_SRAM;
        num_words_cnt_sram <= 0;
        done_cnt_sram <= 0;
        cgra_done_pulse_sram <= 0;
    end
    else if (clk_en) begin
        if (mode == SRAM) begin
            if (cgra_start_pulse) begin
                if ((&num_words) == 1) begin //num_words == {GLB_ADDR_WIDTH{1'b1}}
                    state_sram <= RUN_SRAM_LOOP;
                    num_words_cnt_sram <= num_words;
                    done_cnt_sram <= done_delay;
                    cgra_done_pulse_sram <= 0;
                end
                else if (num_words > 0) begin
                    state_sram <= RUN_SRAM;
                    num_words_cnt_sram <= num_words;
                    done_cnt_sram <= done_delay;
                    cgra_done_pulse_sram <= 0;
                end
                else begin //num_words == 0
                    state_sram <= DONE_SRAM;
                    num_words_cnt_sram <= 0;
                    done_cnt_sram <= done_delay;
                    cgra_done_pulse_sram <= 0;
                end
            end
            else begin
                case (state_sram)
                    IDLE_SRAM: begin
                        state_sram <= IDLE_SRAM;
                        num_words_cnt_sram <= 0;
                        done_cnt_sram <= 0;
                        cgra_done_pulse_sram <= 0;
                    end
                    RUN_SRAM: begin
                        if (cgra_to_io_wr_en_sram == 1 || cgra_to_io_rd_en_sram == 1) begin
                            if (num_words_cnt_sram == 1) begin
                                state_sram <= DONE_SRAM;
                                num_words_cnt_sram <= 0;
                                done_cnt_sram <= done_cnt_sram;
                                cgra_done_pulse_sram <= 0;
                            end
                            else begin
                                state_sram <= RUN_SRAM;
                                num_words_cnt_sram <= num_words_cnt_sram - 1;
                                done_cnt_sram <= done_cnt_sram;
                                cgra_done_pulse_sram <= 0;
                            end
                        end
                        else begin
                            state_sram <= RUN_SRAM;
                            num_words_cnt_sram <= num_words_cnt_sram;
                            done_cnt_sram <= done_cnt_sram;
                            cgra_done_pulse_sram <= 0;
                        end
                    end
                    RUN_SRAM_LOOP: begin
                        state_sram <= RUN_SRAM_LOOP;
                        num_words_cnt_sram <= num_words_cnt_sram;
                        done_cnt_sram <= done_cnt_sram;
                        cgra_done_pulse_sram <= 0;
                    end
                    DONE_SRAM: begin
                        if (done_cnt_sram == 0) begin
                            state_sram <= IDLE_SRAM;
                            num_words_cnt_sram <= 0;
                            done_cnt_sram <= 0;
                            cgra_done_pulse_sram <= 1;
                        end
                        else begin
                            state_sram <= DONE_SRAM;
                            num_words_cnt_sram <= 0;
                            done_cnt_sram <= done_cnt_sram - 1;
                            cgra_done_pulse_sram <= 0;
                        end
                    end
                endcase
            end
        end
        else begin
            state_sram <= IDLE_SRAM;
            num_words_cnt_sram <= 0;
            done_cnt_sram <= 0;
            cgra_done_pulse_sram <= 0;
        end
    end
end

// In SRAM mode, addr comes from cgra with ADDR_OFFSET bits set to 0
assign int_addr_sram = {{cgra_to_io_addr_high[0 +: GLB_ADDR_WIDTH-CGRA_DATA_WIDTH]}, {cgra_to_io_addr_low}};

// We need mux due to the difference BANK_DATA_WIDTH and CGRA_DATA_WIDTH
assign data_sel_sram = int_addr_sram[CGRA_DATA_BYTE-1 +: DATA_SEL_WIDTH];

assign io_to_bank_addr_sram = {int_addr_sram[GLB_ADDR_WIDTH-1:BANK_ADDR_OFFSET], {BANK_ADDR_OFFSET{1'b0}}};
always_comb begin
    if ((state_sram == RUN_SRAM) | (state_sram == RUN_SRAM_LOOP)) begin
        io_to_bank_wr_en_sram = cgra_to_io_wr_en_sram;
        io_to_bank_rd_en_sram = cgra_to_io_rd_en_sram;
        io_to_bank_wr_data_sram = 0;
        io_to_bank_wr_data_sram[data_sel_sram*CGRA_DATA_WIDTH +: CGRA_DATA_WIDTH] = cgra_to_io_wr_data_sram;
        io_to_bank_bit_sel_sram = 0;
        io_to_bank_bit_sel_sram[data_sel_sram*CGRA_DATA_WIDTH +: CGRA_DATA_WIDTH] = {CGRA_DATA_WIDTH{1'b1}};
    end
    else begin
        io_to_bank_rd_en_sram = 0;
        io_to_bank_wr_en_sram = 0;
        io_to_bank_wr_data_sram = 0;
        io_to_bank_bit_sel_sram = 0;
    end
end

// Need mux to select CGRA_DATA from BANK_DATA due to DATA_WIDTH difference
always_ff @(posedge clk) begin
    if (clk_en) begin
        data_sel_sram_d1 <= data_sel_sram;
        data_sel_sram_d2 <= data_sel_sram_d1;
    end
end
assign io_to_cgra_rd_data_sram = int_bank_to_io_rd_data[data_sel_sram_d2 * CGRA_DATA_WIDTH +: CGRA_DATA_WIDTH];

// assign rd_data_valid
always_ff @(posedge clk) begin
    if (clk_en) begin
        io_to_bank_rd_en_sram_d1 <= io_to_bank_rd_en_sram;
        io_to_bank_rd_en_sram_d2 <= io_to_bank_rd_en_sram_d1;
    end
end
assign io_to_cgra_rd_data_valid_sram = int_bank_to_io_rd_data_valid & io_to_bank_rd_en_sram_d2;

//============================================================================//
// output declaration depending on the mode
//============================================================================//
always_comb begin
    case (mode)
        IDLE: begin
            io_to_cgra_rd_data = 0;
            io_to_cgra_rd_data_valid = 0;
            io_to_bank_wr_en = 0;
            io_to_bank_wr_data = 0;
            io_to_bank_wr_data_bit_sel = 0;
            io_to_bank_rd_en = 0;
            io_to_bank_addr = 0;
            cgra_done_pulse = 0;
        end
        INSTREAM: begin
            io_to_cgra_rd_data = io_to_cgra_rd_data_instream;
            io_to_cgra_rd_data_valid = io_to_cgra_rd_data_valid_instream;
            io_to_bank_wr_en = 0;
            io_to_bank_wr_data = 0;
            io_to_bank_wr_data_bit_sel = 0;
            io_to_bank_rd_en = io_to_bank_rd_en_instream;
            io_to_bank_addr = io_to_bank_addr_instream;
            cgra_done_pulse = cgra_done_pulse_instream;
        end
        OUTSTREAM: begin
            io_to_cgra_rd_data = 0;
            io_to_cgra_rd_data_valid = 0;
            io_to_bank_wr_en = io_to_bank_wr_en_outstream;
            io_to_bank_wr_data = io_to_bank_wr_data_outstream;
            io_to_bank_wr_data_bit_sel = io_to_bank_bit_sel_outstream;
            io_to_bank_rd_en = 0;
            io_to_bank_addr = io_to_bank_addr_outstream;
            cgra_done_pulse = cgra_done_pulse_outstream;
        end
        SRAM: begin
            io_to_cgra_rd_data = io_to_cgra_rd_data_sram;
            io_to_cgra_rd_data_valid = io_to_cgra_rd_data_valid_sram;
            io_to_bank_wr_en = io_to_bank_wr_en_sram;
            io_to_bank_wr_data = io_to_bank_wr_data_sram;
            io_to_bank_wr_data_bit_sel = io_to_bank_bit_sel_sram;
            io_to_bank_rd_en = io_to_bank_rd_en_sram;
            io_to_bank_addr = io_to_bank_addr_sram;
            cgra_done_pulse = cgra_done_pulse_sram;
        end
        default: begin
            io_to_cgra_rd_data = 0;
            io_to_cgra_rd_data_valid = 0;
            io_to_bank_wr_en = 0;
            io_to_bank_wr_data = 0;
            io_to_bank_wr_data_bit_sel = 0;
            io_to_bank_rd_en = 0;
            io_to_bank_addr = 0;
            cgra_done_pulse = 0;
        end
    endcase
    if (clk_en == 0) begin
        io_to_bank_wr_en = 0;
        io_to_bank_rd_en = 0;
    end
end

endmodule
