class Config;
    int num_trans;


